/*-----------------------------------------------------------------------------
   Este fichero es parte del procesador DAPA2014 diseñado en la asignatura
   Diseño de Avanzado de Procesadores y Aplicaciones del
   Master Universitario en Ingeniería de Computadores y Redes de la
   Universidad de Sevilla

   It is distributed under GNU General Public License
   See at http://www.gnu.org/licenses/gpl.html
   Copyright (C) 2013 Paulino Ruiz de Clavijo Vázquez <paulino@dte.us.es>
   You can get more info at http://www.dte.us.es/id2
--------------------------------------------------------------------------------

   Fecha:     04-12-2013
   Revisión:  1

   Autor/es:
   Comentarios:

--*--------------------------------- End auto header, don't touch this line --*/
`timescale 1ns / 1ps

module alu(
    input [7:0] a,
    input [7:0] b,
    input [3:0] s_in,
    input [3:0] op,
    output reg s_c,
    output reg s_z,
    output reg s_n,
    output reg s_v,
    output reg [7:0] result
    );

reg[3:0] estado=0;
reg[8:0] tempResult=0;

always @*
	result=tempResult[7:0];

//Modificaci�n de estado
always @* begin
	case (op)
		4'b0000: estado=0;
		4'b0001: estado=1;
		4'b0010: estado=0;
		4'b0011: estado=2;
		4'b0100: estado=3;
		4'b0101: estado=4;
		4'b0110: estado=5;
		4'b0111: estado=5;
		4'b1000: estado=6;
		4'b1001: estado=6;
		4'b1010: estado=7;
		4'b1011: estado=7;
		4'b1100: estado=8;
		4'b1101: estado=8;
		4'b1110: estado=8;
		4'b1111: estado=8;
	endcase
end

//Seg�n el estado
always @* begin
	case (estado)
		0: begin
				tempResult=9'bZZZZZZZZZ;
				s_v=s_in[3];
				s_n=s_in[2];
				s_z=s_in[1];
				s_c=0;
			end
		1: begin
				tempResult=9'bZZZZZZZZZ;
				s_v=1'bZ;
				s_n=1'bZ;
				s_z=1'bZ;
				s_c=1'bZ;
			end
		2: begin
				tempResult=9'bZZZZZZZZZ;
				s_v=s_in[3];
				s_n=s_in[2];
				s_z=s_in[1];
				s_c=1;
			end
		3: begin
				tempResult={1'b0,s_in[0],a[7:1]};  //Sale a[0]
				s_v=s_in[0]^a[0];
				s_n=tempResult[7];
				s_z=((tempResult[7:0]==0)? 1:0);
				s_c=a[0];
			end
		4: begin
				tempResult={1'b0,a[6:0],s_in[0]};  //Sale a[7]
				s_v=a[7]^a[6];
				s_n=tempResult[7];
				s_z=((tempResult[7:0]==0)? 1:0);
				s_c=a[7];
			end
		5: begin
				tempResult=a;
				s_v=1'bZ;
				s_n=1'bZ;
				s_z=1'bZ;
				s_c=1'bZ;
			end
		6: begin  //SUMA
				tempResult=a+b;
				
				//Al sumar dos n�meros complemento dos de distinto signo, el resultado
				//nunca genera un overflow pues la magnitud del n�mero resultante es
				//estrictamente menor que la de cada uno de sus argumentos, y por
				//consiguiente representable. Solo tendremos en cuenta cuando ambos
				//tienen igual signo.
				
				//Al sumar n�meros de igual signo, el overflow se da cuando, como
				//consecuencia de estas rotaciones, el resultado corresponde a un
				//numero de signo contrario al de sus argumentos.
				
				if(a>0 && b>0 && tempResult[7]!=0) //ambos positivos y resultado negativo
					s_v=1;
				else if(a<0 && b<0 && tempResult[7]==0) //ambos negativos y resultado positivo
					s_v=1;
				else
					s_v=0;
				s_n=tempResult[7];
				s_z=((tempResult[7:0]==0)? 1:0);
				s_c=((tempResult[8]==1)? 1:0);
			end
		7: begin  //RESTA
				tempResult=a-b;
				//Underflow:
				if(a>=0 && b<0 && tempResult[7]!=0) //ambos "positivos" (a-b con b neg --> a+b) y resultado negativo
					s_v=1;
				else if(a<=0 && b>0 && tempResult[7]==0) //ambos "negativos" (a-b con a neg y b pos --> -(a+b)) y resultado positivo
					s_v=1;
				else if(a>=0 && b>0 && tempResult[7]!=0) //ambos positivos (a-b con b pos --> a-b) y resultado negativo
					s_v=1;
				else
					s_v=0;
				s_n=tempResult[7];
				s_z=((tempResult[7:0]==0)? 1:0);
				s_c=((tempResult[8]==1)? 1:0);
			end
		8: begin
				tempResult=b;
				s_v=1'bZ;
				s_n=1'bZ;
				s_z=1'bZ;
				s_c=1'bZ;
			end
		default: begin
				tempResult=9'bZZZZZZZZZ;
				s_v=1'bZ;
				s_n=1'bZ;
				s_z=1'bZ;
				s_c=1'bZ;
			end

	endcase
end

endmodule
